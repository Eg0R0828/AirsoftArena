    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   GameManager+DATA   moneyroundsitemsfirst_weaponsecond_weaponstorage  System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   �  �  	      �Base_AK74{PistolGrip_AKPlasticOrange{}Magazine_AK545BunkerPlasticOrange{}Butt_AK74{}Forend_AK74{}ReceiverCover_AKRibbed{}-{}Battery_AKLipo1000{}} 10000 0 0    	      System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	                 	                  