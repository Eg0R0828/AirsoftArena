    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   GameManager+SETTINGS   userNamequalitySettingswindowedMode        Player    